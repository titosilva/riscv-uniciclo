library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.riscv_components.all;

entity RISCV is
  port (
    clock: in std_logic
  );
end RISCV;

architecture RTL of ent is
begin
  --process
end RTL;
