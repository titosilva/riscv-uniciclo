library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

entity ent is
  port (
    --ports
  );
end ent;

architecture RTL of ent is
  --signals
begin
  --process
end RTL;
