library IEEE;
use IEEE.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.riscv_components.all;

entity riscv is
  port (
    clock: in std_logic
  );
end riscv;

architecture RTL of riscv is
begin
  --process
end RTL;
